module mux4_1 (sel, i1, i2, i3, i4, o);
   input [1:0] sel;
   input [15:0] i1, i2, i3, i4;
   output reg [15:0] o;

   always @ (*) begin
      case (sel)
         0: o = i1;
         1: o = i2;
         2: o = i3;
         3: o = i4;
      endcase
   end

endmodule


module mux2_1 (sel, i1, i2, o);
   input sel;
   input [15:0] i1, i2;
   output reg [15:0] o;

   always @ (*) begin
      case (sel)
         0: o = i1;
         1: o = i2;
      endcase
   end

endmodule

module immediate_generator(immediate_value, extended_immediate_value);
    input [7:0] immediate_value;
    output [15:0] extended_immediate_value;
    
    assign extended_immediate_value = {{8{immediate_value[7]}}, immediate_value[7:0]};
endmodule

module counter(clk, reset, on, cnt);
	input clk;
	input reset;
	input on;
	output reg [7:0] cnt;
	always @(*) begin
		if(reset) begin
			cnt = 0;
		end
	end
	always @(posedge clk) begin
		if(on) begin
			cnt <= cnt+ 1;
		end
	end
endmodule